/*Diseña un sistema digital que integre un contador binario de 4 bits y un módulo convertidor binario
a display de 7 segmentos para mostrar el conteo. El sistema debe contar de 0 a 15 con reloj síncrono y
reset asíncrono. El display debe actualizarse con el valor actual del contador. Simula la funcionalidad
completa mostrando señales internas y la salida para el display en GTKWave.*/

module pc_display7s(
    input clk,
    input reset,
    output [6:0] display
  
);

    always

endmodule